
`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////

module adder(
    input [7:0] A_in,
    input [7:0] B_in,
    input Sel_in,
    output [8:0] Rez_out
    );

endmodule
