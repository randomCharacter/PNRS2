`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
module semafor(
    input clk,
    input reset_n,
    input [1:0] Sel_in,
    output [2:0] RGB_A,
    output [2:0] RGB_B
    );


endmodule
